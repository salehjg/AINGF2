-------------------------------------------------------------------------------
--                                                                           --
--          X       X   XXXXXX    XXXXXX    XXXXXX    XXXXXX      X          --
--          XX     XX  X      X  X      X  X      X  X           XX          --
--          X X   X X  X         X      X  X      X  X          X X          --
--          X  X X  X  X         X      X  X      X  X         X  X          --
--          X   X   X  X          XXXXXX   X      X   XXXXXX      X          --
--          X       X  X         X      X  X      X         X     X          --
--          X       X  X         X      X  X      X         X     X          --
--          X       X  X      X  X      X  X      X         X     X          --
--          X       X   XXXXXX    XXXXXX    XXXXXX    XXXXXX      X          --
--                                                                           --
--                                                                           --
--                       O R E G A N O   S Y S T E M S                       --
--                                                                           --
--                            Design & Consulting                            --
--                                                                           --
-------------------------------------------------------------------------------
--                                                                           --
--         Web:           http://www.oregano.at/                             --
--                                                                           --
--         Contact:       mc8051@oregano.at                                  --
--                                                                           --
-------------------------------------------------------------------------------
--                                                                           --
--  MC8051 - VHDL 8051 Microcontroller IP Core                               --
--  Copyright (C) 2001 OREGANO SYSTEMS                                       --
--                                                                           --
--  This library is free software; you can redistribute it and/or            --
--  modify it under the terms of the GNU Lesser General Public               --
--  License as published by the Free Software Foundation; either             --
--  version 2.1 of the License, or (at your option) any later version.       --
--                                                                           --
--  This library is distributed in the hope that it will be useful,          --
--  but WITHOUT ANY WARRANTY; without even the implied warranty of           --
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU        --
--  Lesser General Public License for more details.                          --
--                                                                           --
--  Full details of the license can be found in the file LGPL.TXT.           --
--                                                                           --
--  You should have received a copy of the GNU Lesser General Public         --
--  License along with this library; if not, write to the Free Software      --
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA  --
--                                                                           --
-------------------------------------------------------------------------------
--
--
--         Author:                 Helmut Mayrhofer
--
--         Filename:               mc8051_ram_sim.vhd
--
--         Date of Creation:       Mon Aug  9 12:14:48 1999
--
--         Version:                $Revision: 1.2 $
--
--         Date of Latest Version: $Date: 2002-01-07 12:16:56 $
--
--
--         Description: The mc8051 internal RAM model.
--
--
--
--
-------------------------------------------------------------------------------
architecture sim of mc8051_ram is

   type   ram_type is array (127 downto 0) of unsigned(7 downto 0); 

   signal gpram:        ram_type;             -- general purpose RAM 


begin

------------------------------------------------------------------------------ 
-- ram_read 
------------------------------------------------------------------------------ 
 
  p_read : process (clk, reset)
  begin
    if reset='1' then
      ram_data_o <= "00000000";
    else
      if Rising_Edge(clk) then
        ram_data_o <= std_logic_vector(gpram(conv_integer(unsigned(ram_adr_i))));
      end if;
    end if;
  end process p_read; 

------------------------------------------------------------------------------ 
-- ram_write
------------------------------------------------------------------------------ 

  p_write : process (clk, reset, ram_en_i)
  begin
    if reset='1' then
      gpram <= (others => (others =>'0'));    -- reset every bit
    else
      if Rising_Edge(clk) then
        if ((ram_en_i='1') and (ram_wr_i='1')) then
          gpram(conv_integer(unsigned(ram_adr_i))) <= unsigned(ram_data_i);
        end if;
      end if;
    end if;
  end process p_write;
  
end sim;
